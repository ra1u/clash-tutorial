// Automatically generated Verilog-2001
module SuperLargeNumber_topEntity(input_0
                                 ,output_0);
  input signed [6:0] input_0;
  output [0:0] output_0;
  SuperLargeNumber_topEntity_0 SuperLargeNumber_topEntity_0_inst
  (.eta_i1 (input_0)
  ,.topLet_o (output_0));
endmodule
