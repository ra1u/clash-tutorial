package SuperLargeNumber_types;
  function logic [6:0] signed_7_to_lv(logic signed [6:0] i);
    signed_7_to_lv = i;
  endfunction
  function logic [0:0] logic_vector_1_to_lv(logic [0:0] i);
    logic_vector_1_to_lv = i;
  endfunction
endpackage : SuperLargeNumber_types
